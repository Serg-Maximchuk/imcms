




<!doctype html public "-//W3C//DTD HTML 4.0 Transitional//EN"
"http://www.w3.org/TR/REC-html40/loose.dtd">
<!-- ViewCVS -- http://viewcvs.sourceforge.net/
by Greg Stein -- mailto:gstein@lyra.org -->
<html>
<head>
<title>SourceForge.net CVS Repository - log - cvs: jazzy/jazzy/dict/phonet.sv</title>
<link rel="stylesheet" href="/viewcvs.py/*docroot*/styles.css" type="text/css">
</head>
<body>
<center>
<iframe SRC="http://ads.osdn.com/?op=iframe&position=1&allpositions=1&site_id=2&section=cvs" width="728" height="90" frameborder="0" border="0" MARGINWIDTH="0" MARGINHEIGHT="0" SCROLLING="no"></iframe>
<!-- image audit code -->
<script LANGUAGE="JAVASCRIPT">
<!--
now = new Date();
tail = now.getTime();
document.write("<IMG SRC='http://images-aud.sourceforge.net/pc.gif?l,");
document.write(tail);
document.write("' WIDTH=1 HEIGHT=1 BORDER=0>");
//-->
</SCRIPT>
<noscript>
<img src="http://images-aud.sourceforge.net/pc.gif?l,81677"
WIDTH=1 HEIGHT=1 BORDER=0>
</noscript>
<!-- end audit code -->
</center>
<div class="vc_navheader">
<table width="100%" border="0" cellpadding="0" cellspacing="0">
<tr>
<td align="left"><a href="/viewcvs.py/#dirlist">[cvs]</a> / <a href="/viewcvs.py/jazzy/#dirlist">jazzy</a> / <a href="/viewcvs.py/jazzy/jazzy/#dirlist">jazzy</a> / <a href="/viewcvs.py/jazzy/jazzy/dict/#dirlist">dict</a> / phonet.sv</h1></td>
<td align="right">

&nbsp;

</td>
</tr>
</table>
</div>
<table width="100%">
<tr><td><h1>cvs: jazzy/jazzy/dict/phonet.sv</h1></td>
<td align=right><a href="http://sourceforge.net"><img src="/sourceforge_whitebg.gif" alt="(logo)" border=0 width=136 height=79></a></td></tr>
</table>

<hr noshade>

Default branch: MAIN
<br>
Bookmark a link to HEAD:
(<a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?view=markup">view</a>)
(<a href="/viewcvs.py/*checkout*/jazzy/jazzy/dict/phonet.sv">download</a>)


<br>



 



<hr size=1 noshade>


<a name="rev1.2"></a>
<a name="jEdit_plugin_0-2-1"></a>
<a name="Version_0-5"></a>
<a name="Release-0-5-1"></a>
<a name="Release_0-5"></a>
<a name="version_0-3-0"></a>
<a name="HEAD"></a>


Revision <b>1.2</b>
 -
(<a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?rev=1.2&view=markup">view</a>)
(<a href="/viewcvs.py/*checkout*/jazzy/jazzy/dict/phonet.sv?rev=1.2">download</a>)


(<a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?annotate=1.2">annotate</a>)


- <a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?r1=1.2">[select for diffs]</a>




<br>

<i>Tue Feb  4 21:20:28 2003 UTC</i> (2 years, 10 months ago) by <i>wobban</i>

<br>Branch:

<a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?only_with_tag=MAIN"><b>MAIN</b></a>



<br>CVS Tags:

<a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?only_with_tag=jEdit_plugin_0-2-1"><b>jEdit_plugin_0-2-1</b></a>,

<a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?only_with_tag=Version_0-5"><b>Version_0-5</b></a>,

<a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?only_with_tag=Release-0-5-1"><b>Release-0-5-1</b></a>,

<a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?only_with_tag=Release_0-5"><b>Release_0-5</b></a>,

<a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?only_with_tag=version_0-3-0"><b>version_0-3-0</b></a>,

<a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?only_with_tag=HEAD"><b>HEAD</b></a>






<br>Changes since <b>1.1: +3 -1 lines</b>







<br>Diff to <a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?r1=1.1&amp;r2=1.2">previous 1.1</a>










<pre>Changed to support/use the new GenericSpellDictionary.
</pre>

<hr size=1 noshade>


<a name="rev1.1"></a>
<a name="jEdit_Plugin_0-2-0"></a>


Revision <b>1.1</b>
 -
(<a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?rev=1.1&view=markup">view</a>)
(<a href="/viewcvs.py/*checkout*/jazzy/jazzy/dict/phonet.sv?rev=1.1">download</a>)


(<a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?annotate=1.1">annotate</a>)


- <a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?r1=1.1">[select for diffs]</a>




<br>

<i>Fri Dec 13 22:34:48 2002 UTC</i> (2 years, 11 months ago) by <i>wobban</i>

<br>Branch:

<a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?only_with_tag=MAIN"><b>MAIN</b></a>



<br>CVS Tags:

<a href="/viewcvs.py/jazzy/jazzy/dict/phonet.sv?only_with_tag=jEdit_Plugin_0-2-0"><b>jEdit_Plugin_0-2-0</b></a>















<pre>A Swedish word file and phonetic files for swedish and english. The english is supplied mainly for testing.
</pre>

 



<a name=diff></a>
<hr noshade>
This form allows you to request diffs between any two revisions of
a file. You may select a symbolic revision name using the selection
box or you may type in a numeric name using the type-in text box.
<p>
<form method=get action="/viewcvs.py/jazzy/jazzy/dict/phonet.sv" name=diff_select>

Diffs between
<select name="r1">
<option value="text" selected>Use Text Field</option>

<option value="1.2:version_0-3-0">version_0-3-0</option>

<option value="1.2:jEdit_plugin_0-2-1">jEdit_plugin_0-2-1</option>

<option value="1.1:jEdit_Plugin_0-2-0">jEdit_Plugin_0-2-0</option>

<option value="1.2:Version_0-5">Version_0-5</option>

<option value="1.2:Release_0-5">Release_0-5</option>

<option value="1.2:Release-0-5-1">Release-0-5-1</option>

<option value="1.2:MAIN">MAIN</option>

<option value="1.2:HEAD">HEAD</option>

</select>
<input type="TEXT" size="12" name="tr1" value="1.1"
onChange="document.diff_select.r1.selectedIndex=0">
and
<select name="r2">
<option value="text" selected>Use Text Field</option>

<option value="1.2:version_0-3-0">version_0-3-0</option>

<option value="1.2:jEdit_plugin_0-2-1">jEdit_plugin_0-2-1</option>

<option value="1.1:jEdit_Plugin_0-2-0">jEdit_Plugin_0-2-0</option>

<option value="1.2:Version_0-5">Version_0-5</option>

<option value="1.2:Release_0-5">Release_0-5</option>

<option value="1.2:Release-0-5-1">Release-0-5-1</option>

<option value="1.2:MAIN">MAIN</option>

<option value="1.2:HEAD">HEAD</option>

</select>
<input type="TEXT" size="12" name="tr2" value="1.2"
onChange="document.diff_select.r1.selectedIndex=0">
<br>Type of Diff should be a
<select name="diff_format" onchange="submit()">
<option value="h" selected>Colored Diff</option>
<option value="l" >Long Colored Diff</option>
<option value="u" >Unidiff</option>
<option value="c" >Context Diff</option>
<option value="s" >Side by Side</option>
</select>
<input type=submit value=" Get Diffs "></form>



<hr noshade>
<a name=branch></a>
<form method=GET action="/viewcvs.py/jazzy/jazzy/dict/phonet.sv">

View only Branch:
<select name="only_with_tag" onchange="submit()">
<option value="" selected>Show all branches</option>

<option value="MAIN" >MAIN</option>

</select>
<input type=submit value=" View Branch ">
</form>


<hr noshade>
<a name=logsort></a>
<form method=get action="/viewcvs.py/jazzy/jazzy/dict/phonet.sv">

Sort log by:
<select name="logsort" onchange="submit()">
<option value="cvs" >Not sorted</option>
<option value="date" selected>Commit date</option>
<option value="rev" >Revision</option>
</select>
<input type=submit value=" Sort ">
</form>


<hr noshade>
<table width="100%" border="0" cellpadding="0" cellspacing="0">
<tr>
<td align="left">
<address><a href="http://sourceforge.net/">Back to SourceForge.net</a></address><br />
Powered by <a href="http://viewcvs.sourceforge.net/">ViewCVS 1.0-dev</a>
</td>
<td align="right">
<h3><a target="_blank" href="/viewcvs.py/*docroot*/help_log.html">ViewCVS and CVS Help</a></h3>
</td>
</tr>
</table>
</body>
</html>

